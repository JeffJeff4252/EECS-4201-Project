// ----  Probes  ----
`define PROBE_F_PC f_pc 
`define PROBE_F_INSN f_insn

`define PROBE_D_PC d_pc 
`define PROBE_D_OPCODE d_opcode 
`define PROBE_D_RD d_rd 
`define PROBE_D_FUNCT3 d_funct3 
`define PROBE_D_RS1 d_rs1 
`define PROBE_D_RS2 d_rs2 
`define PROBE_D_FUNCT7 d_funct7 
`define PROBE_D_IMM d_imm 
`define PROBE_D_SHAMT d_imm[4:0]
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd2
// ----  Top module  ----
