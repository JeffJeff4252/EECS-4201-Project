/*
 * Module: decode
 *
 * Description: Decode stage
 *
 * Inputs:
 * 1) clk
 * 2) rst signal
 * 3) insn_iruction ins_i
 * 4) program counter pc_i
 * Outputs:
 * 1) AWIDTH wide program counter pc_o
 * 2) DWIDTH wide insn_iruction output insn_o
 * 3) 5-bit wide destination register ID rd_o
 * 4) 5-bit wide source 1 register ID rs1_o
 * 5) 5-bit wide source 2 register ID rs2_o
 * 6) 7-bit wide funct7 funct7_o
 * 7) 3-bit wide funct3 funct3_o
 * 8) 32-bit wide immediate imm_o
 * 9) 5-bit wide shift amount shamt_o
 * 10) 7-bit width opcode_o
 */

`include "constants.svh"

module decode #(
    parameter int DWIDTH=32,
    parameter int AWIDTH=32
)(
	// inputs
	input logic clk,
	input logic rst,
	input logic [DWIDTH - 1:0] insn_i,
	input logic [DWIDTH - 1:0] pc_i,

    // outputs
    output logic [AWIDTH-1:0] pc_o,
    output logic [DWIDTH-1:0] insn_o,
    output logic [6:0] opcode_o,
    output logic [4:0] rd_o,
    output logic [4:0] rs1_o,
    output logic [4:0] rs2_o,
    output logic [6:0] funct7_o,
    output logic [2:0] funct3_o,
    output logic [4:0] shamt_o,
    output logic [DWIDTH-1:0] imm_o
);

    // Internal signal names (kept as original to preserve top-level naming)
    logic [6:0] opcode, funct7;
    logic [4:0] rs1, rs2, rd, shiftamt;
    logic [2:0] funct3;
    logic [DWIDTH-1:0] instruction, imm_reg;
    logic [AWIDTH-1:0] programcounter;

    // Opcode comes from instruction LSBs
    assign opcode = instruction[6:0];

    // Assign wires for output (drive outputs from local registers)
    assign insn_o = instruction;
    assign pc_o = programcounter;
    assign opcode_o = opcode;
    assign funct3_o = funct3;
    assign funct7_o = funct7;
    assign rs1_o = rs1;
    assign rs2_o = rs2;
    assign rd_o = rd;
    assign shamt_o = shiftamt;

    // Connect inputs to internal registers
    assign instruction = insn_i;
    assign programcounter = pc_i;

    // Combinational decode: extract fields from instruction word
    always_comb begin
        rd = instruction[11:7];
        rs1 = instruction[19:15];
        rs2 = instruction[24:20];
        funct3 = instruction[14:12];
        funct7 = instruction[31:25];
        imm_reg = {{DWIDTH-12{instruction[31]}}, instruction[31:20]};
        shiftamt = instruction[24:20];
    end

endmodule : decode

