/*
 * Module: pd3
 *
 * Description: Top level module that will contain sub-module instantiations.
 *
 * Inputs:
 * 1) clk
 * 2) reset signal
 */


`include "constants.svh"

module pd3 #(
    parameter int AWIDTH = 32,
    parameter int DWIDTH = 32)(
    input logic clk,
    input logic reset
);

    
    // --------------------------------------------------------------------------
    // Control Signals (From Control Unit)
    // --------------------------------------------------------------------------
    logic [DWIDTH-1:0]  CTRL_INSN_I;     // Input instruction for control logic
    logic [6:0]         CTRL_OPCODE_I;   // Opcode extracted from instruction
    logic [6:0]         CTRL_FUNCT7_I;   // Function7 field from instruction
    logic [2:0]         CTRL_FUNCT3_I;   // Function3 field from instruction

    // Control outputs that determine datapath behavior
    logic               CTRL_PCSEL_O;    // Selects next PC (branch or sequential)
    logic               CTRL_IMMSEL_O;   // Selects immediate or register as ALU operand
    logic               CTRL_REGWREN_O;  // Register write enable
    logic               CTRL_RS1SEL_O;   // RS1 selection signal
    logic               CTRL_RS2SEL_O;   // RS2 selection signal
    logic               CTRL_MEMREN_O;   // Memory read enable
    logic               CTRL_MEMWREN_O;  // Memory write enable
    logic [1:0]         CTRL_WBSEL_O;    // Write-back select (e.g., ALU result, memory, etc.)
    logic [3:0]         CTRL_ALUSEL_O;   // ALU operation select

    // --------------------------------------------------------------------------
    // Fetch Stage Signals
    // --------------------------------------------------------------------------
    logic [AWIDTH-1:0]  FETCH_PC_O;      // Program Counter output
    logic [DWIDTH-1:0]  FETCH_INSN_O;    // Instruction fetched from memory

    // --------------------------------------------------------------------------
    // Decode Stage Signals
    // --------------------------------------------------------------------------
    logic [DWIDTH-1:0]  DECODE_INSN_I;   // Input instruction to decode
    logic [AWIDTH-1:0]  DECODE_PC_I;     // Input PC to decode stage

    // Outputs from decode stage
    logic [AWIDTH-1:0]  DECODE_PC_O;
    logic [DWIDTH-1:0]  DECODE_INSN_O;
    logic [6:0]         DECODE_OPCODE_O;
    logic [4:0]         DECODE_RD_O;
    logic [4:0]         DECODE_RS1_O;
    logic [4:0]         DECODE_RS2_O;
    logic [2:0]         DECODE_FUNCT3_O;
    logic [6:0]         DECODE_FUNCT7_O;
    logic [4:0]         DECODE_SHAMT_O;  // Shift amount
    logic [DWIDTH-1:0]  DECODE_IMM_O;    // Immediate value

    // --------------------------------------------------------------------------
    // Immediate Generation (IGEN)
    // --------------------------------------------------------------------------
    logic [6:0]         IGEN_OPCODE_I;
    logic [DWIDTH-1:0]  IGEN_INSN_I;
    logic [DWIDTH-1:0]  IGEN_IMM_O;      // Generated immediate output

    // --------------------------------------------------------------------------
    // Memory Interface
    // --------------------------------------------------------------------------
    logic [AWIDTH-1:0]  MEM_ADDR_I;      // Memory address
    logic [DWIDTH-1:0]  MEM_DATA_I;      // Data input to memory (write data)
    logic               MEM_READ_EN_I;   // Memory read enable
    logic               MEM_WRITE_EN_I;  // Memory write enable
    logic [DWIDTH-1:0]  MEM_DATA_O;      // Memory data output
    logic               MEM_DATA_VLD_O;  // Data valid output

    // --------------------------------------------------------------------------
    // Register File Interface
    // --------------------------------------------------------------------------
    logic [4:0]         RF_RS1_I;        // Register source 1 index
    logic [4:0]         RF_RS2_I;        // Register source 2 index
    logic [4:0]         RF_RD_I;         // Register destination index
    logic [DWIDTH-1:0]  RF_DATAWB_I;     // Data to be written back
    logic               RF_REGWREN_I;    // Register write enable
    logic [DWIDTH-1:0]  RF_RS1DATA_O;    // Output from RS1 register
    logic [DWIDTH-1:0]  RF_RS2DATA_O;    // Output from RS2 register

    // --------------------------------------------------------------------------
    // ALU Interface
    // --------------------------------------------------------------------------
    logic [AWIDTH-1:0]  ALU_PC_I;        // PC input to ALU
    logic [DWIDTH-1:0]  ALU_RS1_I;       // Operand 1
    logic [DWIDTH-1:0]  ALU_RS2_I;       // Operand 2
    logic [3:0]         ALU_SEL_I;       // ALU operation select
    logic [DWIDTH-1:0]  ALU_RES_O;       // ALU result
    logic               ALU_BRTAKEN_O;   // Branch decision

    // --------------------------------------------------------------------------
    // Branch Control Interface
    // --------------------------------------------------------------------------
    logic               BC_OPCODE_I;     // Branch opcode input
    logic               BC_FUNCT3_I;     // Branch funct3 field input
    logic [DWIDTH-1:0]  BC_RS1_I;        // RS1 value for branch comparison
    logic [DWIDTH-1:0]  BC_RS2_I;        // RS2 value for branch comparison
    logic               BC_BREQ_O;       // Branch equal flag
    logic               BC_BRLT_O;       // Branch less-than flag

    // --------------------------------------------------------------------------
    // CONTROL MODULE
    // Generates control signals based on opcode, funct3, funct7, etc.
    // --------------------------------------------------------------------------
    control #(
        .DWIDTH(DWIDTH)
    ) ctrl_inst (
        .insn_i     (CTRL_INSN_I),
        .opcode_i   (CTRL_OPCODE_I),
        .funct7_i   (CTRL_FUNCT7_I),
        .funct3_i   (CTRL_FUNCT3_I),
        .pcsel_o    (CTRL_PCSEL_O),
        .immsel_o   (CTRL_IMMSEL_O),
        .regwren_o  (CTRL_REGWREN_O),
        .rs1sel_o   (CTRL_RS1SEL_O),
        .rs2sel_o   (CTRL_RS2SEL_O),
        .memren_o   (CTRL_MEMREN_O),
        .memwren_o  (CTRL_MEMWREN_O),
        .wbsel_o    (CTRL_WBSEL_O),
        .alusel_o   (CTRL_ALUSEL_O)
    );

    // Control inputs are driven from Decode outputs
    assign CTRL_INSN_I   = DECODE_INSN_O;
    assign CTRL_OPCODE_I = DECODE_OPCODE_O;
    assign CTRL_FUNCT7_I = DECODE_FUNCT7_O;
    assign CTRL_FUNCT3_I = DECODE_FUNCT3_O;

    // --------------------------------------------------------------------------
    // FETCH STAGE
    // Responsible for fetching instructions from memory based on PC.
    // --------------------------------------------------------------------------
    fetch fetch_i(
        .clk    (clk),
        .rst    (reset),
        .pc_o   (FETCH_PC_O),
        .insn_o (FETCH_INSN_O)
    );

    // Fetched instruction comes from memory output
    assign FETCH_INSN_O = MEM_DATA_O;

    // --------------------------------------------------------------------------
    // INSTRUCTION MEMORY
    // Provides instruction words based on PC address.
    // --------------------------------------------------------------------------
    memory #(
        .AWIDTH(AWIDTH),
        .DWIDTH(DWIDTH)
    ) insn_mem (
        .clk        (clk),
        .rst        (reset),
        .addr_i     (MEM_ADDR_I),
        .data_i     (MEM_DATA_I),
        .read_en_i  (MEM_READ_EN_I),
        .write_en_i (MEM_WRITE_EN_I),
        .data_o     (MEM_DATA_O),
        .data_vld_o (MEM_DATA_VLD_O)
    );

    // Memory input signals: always reading instruction memory
    assign MEM_ADDR_I     = DECODE_PC_O;
    assign MEM_DATA_I     = 32'b0;
    assign MEM_READ_EN_I  = 1'b1;
    assign MEM_WRITE_EN_I = 1'b0;

    // --------------------------------------------------------------------------
    // DECODE STAGE
    // Extracts fields such as opcode, rd, rs1, rs2, funct3, funct7, etc.
    // --------------------------------------------------------------------------
    decode decode_i(
        .clk      (clk),
        .rst      (reset),
        .insn_i   (DECODE_INSN_I),
        .pc_i     (DECODE_PC_I),
        .pc_o     (DECODE_PC_O),
        .insn_o   (DECODE_INSN_O),
        .opcode_o (DECODE_OPCODE_O),
        .rd_o     (DECODE_RD_O),
        .rs1_o    (DECODE_RS1_O),
        .rs2_o    (DECODE_RS2_O),
        .funct3_o (DECODE_FUNCT3_O),
        .funct7_o (DECODE_FUNCT7_O),
        .shamt_o  (DECODE_SHAMT_O),
        .imm_o    (DECODE_IMM_O)
    );

    assign DECODE_INSN_I = FETCH_INSN_O;
    assign DECODE_PC_I   = FETCH_PC_O;
    assign DECODE_IMM_O  = IGEN_IMM_O;

    // --------------------------------------------------------------------------
    // IMMEDIATE GENERATOR (IGEN)
    // Extracts and formats immediates depending on instruction type.
    // --------------------------------------------------------------------------
    igen igen_i(
        .opcode_i (IGEN_OPCODE_I),
        .insn_i   (IGEN_INSN_I),
        .imm_o    (IGEN_IMM_O)
    );

    assign IGEN_OPCODE_I = DECODE_OPCODE_O;
    assign IGEN_INSN_I   = DECODE_INSN_O;

    // --------------------------------------------------------------------------
    // REGISTER FILE
    // Holds 32 general-purpose registers.
    // Provides two read ports and one write port.
    // --------------------------------------------------------------------------
    register_file #(
        .DWIDTH(DWIDTH)
    ) register_file_i (
        .clk        (clk),
        .rst        (reset),
        .rs1_i      (RF_RS1_I),
        .rs2_i      (RF_RS2_I),
        .rd_i       (RF_RD_I),
        .datawb_i   (RF_DATAWB_I),
        .regwren_i  (RF_REGWREN_I),
        .rs1data_o  (RF_RS1DATA_O),
        .rs2data_o  (RF_RS2DATA_O)
    );

    assign RF_RS1_I     = DECODE_RS1_O;
    assign RF_RS2_I     = DECODE_RS2_O;
    assign RF_RD_I      = DECODE_RD_O;
    assign RF_DATAWB_I  = 'd0;                // No writeback yet connected
    assign RF_REGWREN_I = CTRL_REGWREN_O;

    // --------------------------------------------------------------------------
    // BRANCH CONTROL
    // Handles comparison logic for branch instructions.
    // Outputs flags for equality and less-than conditions.
    // --------------------------------------------------------------------------
    branch_control branching(
        .opcode_i (DECODE_OPCODE_O),
        .funct3_i (DECODE_FUNCT3_O),
        .rs1_i    (RF_RS1DATA_O),
        .rs2_i    (RF_RS2DATA_O),
        .breq_o   (BC_BREQ_O),
        .brlt_o   (BC_BRLT_O)
    );

    assign BC_OPCODE_I = DECODE_OPCODE_O;
    assign BC_FUNCT3_I = DECODE_FUNCT3_O;
    assign BC_RS1_I    = RF_RS1DATA_O;
    assign BC_RS2_I    = RF_RS2DATA_O;

    // --------------------------------------------------------------------------
    // BRANCH DECISION LOGIC
    // Determines whether to take a branch based on instruction type and condition flags.
    // --------------------------------------------------------------------------
    always_comb begin : BRANCHER
        if (DECODE_OPCODE_O == BRANCH) begin
            case (DECODE_FUNCT3_O)
                'h0: ALU_BRTAKEN_O = BC_BREQ_O;       // BEQ
                'h1: ALU_BRTAKEN_O = ~BC_BREQ_O;      // BNE
                'h4, 'h6: ALU_BRTAKEN_O = BC_BRLT_O;  // BLT / BLTU
                'h5, 'h7: ALU_BRTAKEN_O = ~BC_BRLT_O; // BGE / BGEU
                default: ALU_BRTAKEN_O = 'd0;
            endcase
        end else begin
            ALU_BRTAKEN_O = 'd0;
        end
    end

    // --------------------------------------------------------------------------
    // ALU
    // Performs arithmetic, logical, and comparison operations.
    // --------------------------------------------------------------------------
    alu #(
        .DWIDTH(DWIDTH),
        .AWIDTH(AWIDTH)
    ) alu_e (
        .pc_i      (ALU_PC_I),
        .funct3_i  (DECODE_FUNCT3_O),
        .funct7_i  (DECODE_FUNCT7_O),
        .rs1_i     (ALU_RS1_I),
        .rs2_i     (ALU_RS2_I),
        .alusel_i  (ALU_SEL_I),
        .res_o     (ALU_RES_O),
        .brtaken_o (ALU_BRTAKEN_O)
    );

    // ALU input selection logic
    assign ALU_PC_I  = DECODE_PC_O;
    assign ALU_RS1_I = RF_RS1DATA_O;
    assign ALU_RS2_I = (CTRL_IMMSEL_O) ? IGEN_IMM_O : RF_RS2DATA_O;
    assign ALU_SEL_I = CTRL_ALUSEL_O;

endmodule : pd3
